library verilog;
use verilog.vl_types.all;
entity stopwatch_vlg_check_tst is
    port(
        clk_out         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end stopwatch_vlg_check_tst;
