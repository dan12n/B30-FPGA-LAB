library verilog;
use verilog.vl_types.all;
entity stopwatchtimes_vlg_vec_tst is
end stopwatchtimes_vlg_vec_tst;
