library verilog;
use verilog.vl_types.all;
entity registeredmultiplier_vlg_vec_tst is
end registeredmultiplier_vlg_vec_tst;
