library verilog;
use verilog.vl_types.all;
entity stopwatch_vlg_vec_tst is
end stopwatch_vlg_vec_tst;
